module adder(
    input  logic a, b, cin,
    output logic sum, cout
);

always_comb begin
    sum  = a ^ b ^ cin;
    cout = (a & b) | (cin & (a ^ b));
end

endmodule
