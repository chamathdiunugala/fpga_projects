`timescale 1ns/1ps

module adder_tb;

    // Testbench signals
    reg a, b, cin;
    reg sum, cout;

    // Instantiate the DUT (Device Under Test)
    adder dut (
        .a(a),
        .b(b),
        .cin(cin),
        .sum(sum),
        .cout(cout)
    );

    // Apply all possible input combinations
    initial begin
        $display("a b cin | sum cout");
        $display("------------------");

        for (int i = 0; i < 8; i++) begin
            {a, b, cin} = i;
            #1; // small delay for propagation
            $display("%b %b  %b  |  %b   %b", a, b, cin, sum, cout);
        end

        $finish;
    end

endmodule
